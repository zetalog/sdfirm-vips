//
// Copyright (c) 1999-2000 Pinhas Krengel.  Permission to copy is granted
// provided that this header remains intact.  This software is provided
// with no warranties.
//

`include "TimeScale.v"
//4096 x 4 ROM + sample + shift and enable logic
module sd_slv_rom(a, e, s, q, ck);
  input  [ 9:0] a; //address
  input         e; //enable
  input         s; //shift
  output [ 3:0] q;
  input         ck;

  wire   [15:0] O;
  wire   [ 3:0] d;
  reg    [ 3:0] q;

  // synthesis translate_off
  initial q=4'hf;
  // synthesis translate_on
  always @ (posedge ck) q <= d;
  
  assign d=
  (e && ~s && a[9:8] == 2'h0) ? O[ 3: 0] :
  (e && ~s && a[9:8] == 2'h1) ? O[ 7: 4] :
  (e && ~s && a[9:8] == 2'h2) ? O[11: 8] :
  (e && ~s && a[9:8] == 2'h3) ? O[15:12] :
  (e &&  s                  ) ? {q[0], q[3:1]} : 
  4'b1111; //drive 0 in order to start with start bit of 0.
                     
  
  defparam u_rom0.INIT=
  256'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010;
  defparam u_rom1.INIT=
  256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001101;
  defparam u_rom2.INIT=
  256'b1111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000;
  defparam u_rom3.INIT=
  256'b1111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000001;
  defparam u_rom4.INIT=
  256'b1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000;
  defparam u_rom5.INIT=
  256'b1111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000;
  defparam u_rom6.INIT=
  256'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
  defparam u_rom7.INIT=
  256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //
  defparam u_rom8.INIT=
  256'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010;
  defparam u_rom9.INIT=
  256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
  defparam u_rom10.INIT=
  256'b1111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000;
  defparam u_rom11.INIT=
  256'b1111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000;
  defparam u_rom12.INIT=
  256'b1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000;
  defparam u_rom13.INIT=
  256'b1111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000;
  defparam u_rom14.INIT=
  256'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
  defparam u_rom15.INIT=
  256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  //
  ROM256X1 u_rom0 (
   .O (O[0]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom0
  ROM256X1 u_rom1 (
   .O (O[1]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom1
  ROM256X1 u_rom2 (
   .O (O[2]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom2
  ROM256X1 u_rom3 (
   .O (O[3]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom3
  ROM256X1 u_rom4 (
   .O (O[4]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom4
  ROM256X1 u_rom5 (
   .O (O[5]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom5
  ROM256X1 u_rom6 (
   .O (O[6]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom6
  ROM256X1 u_rom7 (
   .O (O[7]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom7
  ROM256X1 u_rom8 (
   .O (O[8]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom8
  ROM256X1 u_rom9 (
   .O (O[9]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom9
  ROM256X1 u_rom10 (
   .O (O[10]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom10
  ROM256X1 u_rom11 (
   .O (O[11]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom11
  ROM256X1 u_rom12 (
   .O (O[12]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom12
  ROM256X1 u_rom13 (
   .O (O[13]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom13
  ROM256X1 u_rom14 (
   .O (O[14]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom14
  ROM256X1 u_rom15 (
   .O (O[15]),
   .A0(a[0]), 
   .A1(a[1]), 
   .A2(a[2]), 
   .A3(a[3]), 
   .A4(a[4]), 
   .A5(a[5]), 
   .A6(a[6]), 
   .A7(a[7])
  );//ROM256X1 u_rom15

endmodule

